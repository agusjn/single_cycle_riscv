//pc_sel = 0 -> chÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â»ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Ân PC + 4 ngÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â°ÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â»ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â£c lÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚ÂºÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡i chÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â»ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Ân PC + IMME
//opa_sel = 0 -> chÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â»ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Ân PC ngÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â°ÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â»ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â£c lÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚ÂºÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡i chÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â»ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Ân rs1
//opb_sel = 0 -> chÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â»ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Ân rs2 ngÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â°ÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â»ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â£c lÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚ÂºÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡i chÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â»ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Ân IMME
//br_un = 0 -> signed ngÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â°ÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â»ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â£c lÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚ÂºÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡i unsigned
//rd_wren = 0 -> khÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â´ng store vÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â o rd ngÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â°ÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â»ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â£c lÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚ÂºÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡i store vÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â o rd
//mem_wren = 0 -> khÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â´ng store vÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â o LSU ngÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â°ÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â»ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â£c lÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚ÂºÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡i store vÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â o LSU
//mem_us = 0 -> signed ngÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â°ÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â»ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â£c lÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚ÂºÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡i unsigned
//wb_sel = 0 -> pc_four, = 1 -> alu data, = 2 -> lsu data



module unit(
    input logic [31:0] instr,
    input logic br_less, 
	 input logic br_equal,
	 
    output logic pc_sel, 
	 output logic opa_sel, 
	 output logic opb_sel, 
	 output logic br_un, 
	 output logic insn_vld, 
	 output logic rd_wren, 
	 output logic mem_wren, 
	 output logic mem_us,
    output logic [3:0] alu_op, 
	 output logic [3:0] mem_wrnum,
    output logic [1:0] wb_sel

    );

 localparam  OP_LOAD  = 7'b00000_11;  // load opcode
 localparam  OP_ALU_I = 7'b00100_11;  // i-type alu opcode
 localparam  OP_AUIPC = 7'b00101_11;  // add upper immediate to pc
 localparam  OP_STORE = 7'b01000_11;  // store opcode
 localparam  OP_ALU_R = 7'b01100_11;  // r-type alu opcode
 localparam  OP_LUI   = 7'b01101_11;  // load upper immediate
 localparam  OP_BR    = 7'b11000_11;  // brach opcode
 localparam  OP_JALR  = 7'b11001_11;  // jump and link reg
 localparam  OP_JAL   = 7'b11011_11;  // jump and link
localparam BEQ = 3'b000;
localparam BNE = 3'b001;
localparam BLT = 3'b100;
localparam BGE = 3'b101;
localparam BLTU = 3'b110;
localparam BGEU = 3'b111;

localparam  LB  = 3'b000;
localparam  LH  = 3'b001;
localparam  LW  = 3'b010;
localparam  LBU = 3'b100;
localparam  LHU = 3'b101;

localparam  SB = 3'b000;
localparam  SH = 3'b001;
localparam  SW = 3'b010;

logic [6:0] opcode ;
logic [2:0] funct3 ;
logic funct7 ;

assign    funct3 = instr[14:12];
assign   funct7 = instr[30];
assign    opcode = instr[6:0];  


always_comb begin 
    case(opcode) 
        OP_ALU_R: begin  //R-type
                pc_sel = 1'b0;
                rd_wren = 1'b1;
                opa_sel = 1'b1;  
                opb_sel = 1'b0;
                wb_sel = 2'd1; //data from ALU
                mem_wren = 1'b0;
                mem_wrnum = 4'b0000;
                mem_us = 1'bx;
                br_un = 1'bx;
                insn_vld = 1'b1;
                case(funct3)
               3'b000: alu_op = (funct7) ? 4'd1 : 4'd0;
               3'b001:	alu_op = 4'd7;
					3'b010:	alu_op = 4'd2;
					3'b011:	alu_op = 4'd3;
					3'b100:	alu_op = 4'd4;
					3'b101: alu_op = (funct7) ? 4'd9 : 4'd8;
					3'b110:	alu_op = 4'd5;
					3'b111:	alu_op = 4'd6;
                    default: alu_op = 4'bxxxx;
                endcase

        end
        OP_ALU_I: begin //I-TYPE
            pc_sel = 1'b0;
            rd_wren = 1'b1;
            opb_sel = 1'b1;
            opa_sel = 1'b1;
            wb_sel = 2'd1;
            mem_wren = 1'b0;
            mem_wrnum = 4'b0000;
            mem_us = 1'bx;
            br_un = 1'bx;
            insn_vld = 1'b1;
            case(funct3)
            3'b000: alu_op = 4'd0;    //addi
				3'b010:	alu_op = 4'd2;    //slti
				3'b011:	alu_op = 4'd3;    //sltiu
				3'b100:	alu_op = 4'd4;    //xori
				3'b110: alu_op = 4'd5;    //ori
				3'b111:	alu_op = 4'd6;    //andi
				3'b001:	alu_op = 4'd7;    //slli
            3'b101: alu_op = (funct7) ? 4'd9 : 4'd8;
                default: alu_op = 4'bxxxx;
            endcase
        end

        7'b0000011: begin //LOAD INSTRUCTION
            pc_sel = 1'b0;
            mem_wren = 1'b0; // not store
            br_un = 1'bx;
            rd_wren = 1'b1;   //write to rd
            opa_sel = 1'b1;   //RS1
            opb_sel = 1'b1;   //IMME
            alu_op = 4'd0;    //add
            wb_sel = 2'd2;    //writeback LSU
             case ( funct3 )
                    LB :    begin
                                mem_wrnum   = 4'b0001; // byte
                                mem_us     = 1'b0;    // sign_ext
                                insn_vld = 1'b1;
                            end
                    LH :    begin
                                mem_wrnum   = 4'b0011; // half-word
                                mem_us   = 1'b0;    // sign_ext
                                insn_vld = 1'b1;
                            end
                    LW :    begin
                                mem_wrnum  = 4'b1111; // word
                                mem_us  = 1'b0;    // sign_ext
                                insn_vld = 1'b1;
                            end
                    LBU:    begin
                                mem_wrnum = 4'b0001; // byte
                                mem_us = 1'b1;    // zero_ext
                                insn_vld = 1'b1;
                            end  
                    LHU:    begin
                                mem_wrnum = 4'b0011; // half-word
                                mem_us = 1'b1;    // zero_ext
                                insn_vld = 1'b1;
                            end
                    default:begin
                                mem_wrnum  = 4'b0;
                                mem_us  = 1'b0;
                                insn_vld = 1'b0;
                             end
            endcase
        end


        OP_STORE: begin //S-TYPE instructions
            pc_sel =1'b0;
            wb_sel = 2'd1;
            mem_us = 1'bx;
            br_un = 1'bx;
            mem_wren = 1'b1; //WRITE LSU
            alu_op = 4'd0;    //add
            rd_wren = 1'b0; // NO Write back
            opa_sel = 1'b1;   //RS1
            opb_sel = 1'b1; //IMME
            case ( funct3 )
                    SB :    begin
                            mem_wrnum   = 4'b0001; // byte
                            insn_vld = 1'b1;
                    end
                    SH :    begin
                            mem_wrnum   = 4'b0011; // half-word
                            insn_vld = 1'b1;
                    end
                    SW :    begin
                            mem_wrnum   = 4'b1111; // word
                            insn_vld = 1'b1;
                    end
                    default: begin
                            mem_wrnum = 4'b0000;
                             insn_vld = 1'b0;
                    end
            endcase
        end



        OP_BR: begin	// B-type instructions
            mem_wren = 1'b0;  //READ MEM
            rd_wren = 1'b0;   //no writeback
            alu_op = 1'b0;    //ADD
            mem_wrnum = 4'b0000;
            mem_us = 1'bx;
				wb_sel = 2'd1;
            opa_sel = 1'b0; //PC
            opb_sel = 1'b1; //IMM
            case(funct3)
            BEQ: begin //beq
                    insn_vld = 1'b1;
                    br_un = 1'b0;
                    pc_sel = (br_equal) ? 1'b1 : 1'b0;
            end
            BNE: begin   //bne
                    insn_vld = 1'b1;
                    br_un = 1'b0;
                    pc_sel = (!br_equal) ? 1'b1 : 1'b0;
            end
            BLT: begin   //blt
                    br_un = 1'b0;
                    insn_vld = 1'b1;
                    pc_sel = (br_less) ? 1'b1 : 1'b0;
            end
            BGE: begin   //bge
                    br_un = 1'b0;
                    insn_vld = 1'b1;
                    pc_sel = ((!br_less && !br_equal ) || br_equal) ? 1'b1 : 1'b0;
            end 
            BLTU: begin   //bltu
                    br_un = 1'b1;
                    insn_vld = 1'b1;
                    pc_sel = (br_less) ? 1'b1 : 1'b0;
            end
            BGEU: begin   //bgeu
                    insn_vld = 1'b1;
                    br_un = 1'b1;
                    pc_sel = ((!br_less && !br_equal ) || br_equal) ? 1'b1 : 1'b0;
            end 
            default:begin
                    br_un = 1'bx;
                    pc_sel = 1'bx;
                    insn_vld = 1'b0;
            end
            endcase
            
        end


        OP_AUIPC: begin	// AUIPC
            insn_vld = 1'b1;
    		rd_wren = 1'b1;
    		opa_sel = 1'b0;       //PC
    		opb_sel = 1'b1;   //IMM
    		mem_wren = 1'b0;  //READ
    		wb_sel = 2'd1;    //ALU
    		alu_op = 4'd0;    //ADD
            pc_sel = 1'b0; //PC+4   
            mem_wrnum = 4'b0000;
            mem_us = 1'bx;
            br_un = 1'bx;
        end
        OP_LUI : begin //LUI
            insn_vld = 1'b1;
            pc_sel = 1'b0;  //PC +4
            rd_wren = 1'b1;   //write
            opa_sel = 1'bx;
            opb_sel = 1'b1; //IMME
            alu_op = 4'd0;
            mem_wren = 1'b0; //not store 
            wb_sel = 2'd1; //ALU
            mem_wrnum = 4'b0000;
            mem_us = 1'bx;
            br_un = 1'bx;
        end
		OP_JAL: begin	// JAL
            insn_vld = 1'b1;
            rd_wren = 1'b1;   
    		opa_sel = 1'b0;   //PC
    		opb_sel = 1'b1;   //IMME
            alu_op = 4'd0;    //ADD
            mem_wren = 1'b0;  // READ
            wb_sel = 2'd0;  //PC + 4 luu vao regfile
            pc_sel = 1'b1; // PC + IMME
            mem_wrnum = 4'bxxxx;
            mem_us = 1'bx;
            br_un = 1'bx;
    		end    
        
        OP_JALR: begin   //JALR
            insn_vld = 1'b1;
            rd_wren = 1'b1;   
    		opa_sel = 1'b1;   //RS1
    		opb_sel = 1'b1;   //IMME
            alu_op = 4'd0;    //ADD
            mem_wren = 1'b0;  // READ
            wb_sel = 2'd0;  //PC + 4 luu vao regfile
            pc_sel = 1'b1; // PC + IMME
            mem_wrnum = 4'bxxxx;
            mem_us = 1'bx;
            br_un = 1'bx;
        end    
        default:  begin 
            insn_vld = 1'b0;         
            rd_wren = 1'b0;   
				opa_sel = 1'b0;   //RS1
				opb_sel = 1'b0;   //IMME
            alu_op = 4'b0;    //ADD
            mem_wren = 1'b0;  // READ
            wb_sel = 2'bxx;  //PC + 4 luu vao regfile
            pc_sel = 1'b0; // PC + IMME
            mem_wrnum = 4'b000;
            mem_us = 1'b0;
            br_un = 1'b0;
        end
    endcase
end


endmodule